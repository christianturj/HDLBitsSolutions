module top_module(
    input clk,
    input in,
    input areset,
    output out); //
    reg[1:0] state, next_state;
    parameter [1:0] A=2'd0; 
    parameter [1:0]B=2'd1; 
    parameter [1:0]C=2'd2;
    parameter [1:0]D=2'd3;
    // State transition logic
    always @ (*)
        begin
            case(state)
                A: next_state=(in ? B : A);
                B: next_state=(in ? B: C);
                C: next_state=(in ? D : A);
                D: next_state=(in ? B: C);
                default: next_state=A;
            endcase
        end
    // State flip-flops with asynchronous reset
    always @(posedge clk or posedge areset)
                begin
                    if(areset)
                        begin
                            state<=A;
                        end
                    else
                        begin
                            state<=next_state;
                        end
                end
                    
    // Output logic
    assign out=(state==D);

endmodule
